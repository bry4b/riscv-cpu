module reorder_buffer #(
    parameter ROB_SIZE = 16,
    parameter COMMIT_PORTS = 1
) (

);

endmodule