module issue_queue #(
    parameter IQ_SIZE = 16,
    parameter ISSUE_PORTS = 2,
    parameter INSTR_SIZE = 32
) (

);


endmodule