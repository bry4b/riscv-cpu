`ifndef _parameters_svh
`define _parameters_svh

parameter NUM_REG = 32;
parameter REG_SIZE = $clog2(NUM_REG);
parameter INSTR_SIZE = 32;

`endif
