module issue_select (

);

endmodule