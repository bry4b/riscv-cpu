module loadstore_queue #(
    parameter LSQ_SIZE = 16,
    parameter INSTR_SIZE = 32
) (

);

endmodule