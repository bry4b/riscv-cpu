`ifndef _parameters_svh
`define _parameters_svh

parameter INSTR_SIZE = 32;

`endif
