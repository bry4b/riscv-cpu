module arch_regfile #(
    parameter NUM_REG = 32,
    parameter REG_SIZE = 32
) (

);

endmodule